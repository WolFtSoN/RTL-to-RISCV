/*
Simple memory-mapped interface

Simple memory model (e.g., small memory array)
*/