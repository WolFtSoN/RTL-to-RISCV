import all_pkgs::*;

module id_ex (
    input logic             id_pc,
    input logic [WIDTH-1:0] reg_data1, reg_data2,
    input logic [WIDTH-1:0] imm_ext
);
    
endmodule