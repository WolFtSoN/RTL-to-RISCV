package a01_defines_pkg;

parameter ADDR_W = 32;
parameter DATA_W = 32;
parameter FIFO_DEPTH = 16;
parameter FIFO_DATA_W = 65;
    
endpackage