/*
Connects everything together
*/